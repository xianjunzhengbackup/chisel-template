module FileReader(
  input        clock,
  input        reset,
  input  [7:0] io_address,
  output [7:0] io_data
);
  wire [7:0] _GEN_1 = 8'h1 == io_address ? 8'h1 : 8'h0; // @[FileReader.scala 21:{11,11}]
  wire [7:0] _GEN_2 = 8'h2 == io_address ? 8'h2 : _GEN_1; // @[FileReader.scala 21:{11,11}]
  wire [7:0] _GEN_3 = 8'h3 == io_address ? 8'h3 : _GEN_2; // @[FileReader.scala 21:{11,11}]
  wire [7:0] _GEN_4 = 8'h4 == io_address ? 8'h4 : _GEN_3; // @[FileReader.scala 21:{11,11}]
  wire [7:0] _GEN_5 = 8'h5 == io_address ? 8'h5 : _GEN_4; // @[FileReader.scala 21:{11,11}]
  wire [7:0] _GEN_6 = 8'h6 == io_address ? 8'h6 : _GEN_5; // @[FileReader.scala 21:{11,11}]
  wire [7:0] _GEN_7 = 8'h7 == io_address ? 8'h7 : _GEN_6; // @[FileReader.scala 21:{11,11}]
  wire [7:0] _GEN_8 = 8'h8 == io_address ? 8'h8 : _GEN_7; // @[FileReader.scala 21:{11,11}]
  wire [7:0] _GEN_9 = 8'h9 == io_address ? 8'h9 : _GEN_8; // @[FileReader.scala 21:{11,11}]
  wire [7:0] _GEN_10 = 8'ha == io_address ? 8'ha : _GEN_9; // @[FileReader.scala 21:{11,11}]
  wire [7:0] _GEN_11 = 8'hb == io_address ? 8'hb : _GEN_10; // @[FileReader.scala 21:{11,11}]
  wire [7:0] _GEN_12 = 8'hc == io_address ? 8'hc : _GEN_11; // @[FileReader.scala 21:{11,11}]
  wire [7:0] _GEN_13 = 8'hd == io_address ? 8'hd : _GEN_12; // @[FileReader.scala 21:{11,11}]
  wire [7:0] _GEN_14 = 8'he == io_address ? 8'he : _GEN_13; // @[FileReader.scala 21:{11,11}]
  wire [7:0] _GEN_15 = 8'hf == io_address ? 8'hf : _GEN_14; // @[FileReader.scala 21:{11,11}]
  wire [7:0] _GEN_16 = 8'h10 == io_address ? 8'h10 : _GEN_15; // @[FileReader.scala 21:{11,11}]
  wire [7:0] _GEN_17 = 8'h11 == io_address ? 8'h11 : _GEN_16; // @[FileReader.scala 21:{11,11}]
  wire [7:0] _GEN_18 = 8'h12 == io_address ? 8'h12 : _GEN_17; // @[FileReader.scala 21:{11,11}]
  wire [7:0] _GEN_19 = 8'h13 == io_address ? 8'h13 : _GEN_18; // @[FileReader.scala 21:{11,11}]
  wire [7:0] _GEN_20 = 8'h14 == io_address ? 8'h14 : _GEN_19; // @[FileReader.scala 21:{11,11}]
  wire [7:0] _GEN_21 = 8'h15 == io_address ? 8'h15 : _GEN_20; // @[FileReader.scala 21:{11,11}]
  wire [7:0] _GEN_22 = 8'h16 == io_address ? 8'h16 : _GEN_21; // @[FileReader.scala 21:{11,11}]
  wire [7:0] _GEN_23 = 8'h17 == io_address ? 8'h17 : _GEN_22; // @[FileReader.scala 21:{11,11}]
  wire [7:0] _GEN_24 = 8'h18 == io_address ? 8'h18 : _GEN_23; // @[FileReader.scala 21:{11,11}]
  wire [7:0] _GEN_25 = 8'h19 == io_address ? 8'h19 : _GEN_24; // @[FileReader.scala 21:{11,11}]
  wire [7:0] _GEN_26 = 8'h1a == io_address ? 8'h1a : _GEN_25; // @[FileReader.scala 21:{11,11}]
  wire [7:0] _GEN_27 = 8'h1b == io_address ? 8'h1b : _GEN_26; // @[FileReader.scala 21:{11,11}]
  wire [7:0] _GEN_28 = 8'h1c == io_address ? 8'h1c : _GEN_27; // @[FileReader.scala 21:{11,11}]
  wire [7:0] _GEN_29 = 8'h1d == io_address ? 8'h1d : _GEN_28; // @[FileReader.scala 21:{11,11}]
  wire [7:0] _GEN_30 = 8'h1e == io_address ? 8'h1e : _GEN_29; // @[FileReader.scala 21:{11,11}]
  wire [7:0] _GEN_31 = 8'h1f == io_address ? 8'h1f : _GEN_30; // @[FileReader.scala 21:{11,11}]
  wire [7:0] _GEN_32 = 8'h20 == io_address ? 8'h20 : _GEN_31; // @[FileReader.scala 21:{11,11}]
  wire [7:0] _GEN_33 = 8'h21 == io_address ? 8'h21 : _GEN_32; // @[FileReader.scala 21:{11,11}]
  wire [7:0] _GEN_34 = 8'h22 == io_address ? 8'h22 : _GEN_33; // @[FileReader.scala 21:{11,11}]
  wire [7:0] _GEN_35 = 8'h23 == io_address ? 8'h23 : _GEN_34; // @[FileReader.scala 21:{11,11}]
  wire [7:0] _GEN_36 = 8'h24 == io_address ? 8'h24 : _GEN_35; // @[FileReader.scala 21:{11,11}]
  wire [7:0] _GEN_37 = 8'h25 == io_address ? 8'h25 : _GEN_36; // @[FileReader.scala 21:{11,11}]
  wire [7:0] _GEN_38 = 8'h26 == io_address ? 8'h26 : _GEN_37; // @[FileReader.scala 21:{11,11}]
  wire [7:0] _GEN_39 = 8'h27 == io_address ? 8'h27 : _GEN_38; // @[FileReader.scala 21:{11,11}]
  wire [7:0] _GEN_40 = 8'h28 == io_address ? 8'h28 : _GEN_39; // @[FileReader.scala 21:{11,11}]
  wire [7:0] _GEN_41 = 8'h29 == io_address ? 8'h29 : _GEN_40; // @[FileReader.scala 21:{11,11}]
  wire [7:0] _GEN_42 = 8'h2a == io_address ? 8'h2a : _GEN_41; // @[FileReader.scala 21:{11,11}]
  wire [7:0] _GEN_43 = 8'h2b == io_address ? 8'h2b : _GEN_42; // @[FileReader.scala 21:{11,11}]
  wire [7:0] _GEN_44 = 8'h2c == io_address ? 8'h2c : _GEN_43; // @[FileReader.scala 21:{11,11}]
  wire [7:0] _GEN_45 = 8'h2d == io_address ? 8'h2d : _GEN_44; // @[FileReader.scala 21:{11,11}]
  wire [7:0] _GEN_46 = 8'h2e == io_address ? 8'h2e : _GEN_45; // @[FileReader.scala 21:{11,11}]
  wire [7:0] _GEN_47 = 8'h2f == io_address ? 8'h2f : _GEN_46; // @[FileReader.scala 21:{11,11}]
  wire [7:0] _GEN_48 = 8'h30 == io_address ? 8'h30 : _GEN_47; // @[FileReader.scala 21:{11,11}]
  wire [7:0] _GEN_49 = 8'h31 == io_address ? 8'h31 : _GEN_48; // @[FileReader.scala 21:{11,11}]
  wire [7:0] _GEN_50 = 8'h32 == io_address ? 8'h32 : _GEN_49; // @[FileReader.scala 21:{11,11}]
  wire [7:0] _GEN_51 = 8'h33 == io_address ? 8'h33 : _GEN_50; // @[FileReader.scala 21:{11,11}]
  wire [7:0] _GEN_52 = 8'h34 == io_address ? 8'h34 : _GEN_51; // @[FileReader.scala 21:{11,11}]
  wire [7:0] _GEN_53 = 8'h35 == io_address ? 8'h35 : _GEN_52; // @[FileReader.scala 21:{11,11}]
  wire [7:0] _GEN_54 = 8'h36 == io_address ? 8'h36 : _GEN_53; // @[FileReader.scala 21:{11,11}]
  wire [7:0] _GEN_55 = 8'h37 == io_address ? 8'h37 : _GEN_54; // @[FileReader.scala 21:{11,11}]
  wire [7:0] _GEN_56 = 8'h38 == io_address ? 8'h38 : _GEN_55; // @[FileReader.scala 21:{11,11}]
  wire [7:0] _GEN_57 = 8'h39 == io_address ? 8'h39 : _GEN_56; // @[FileReader.scala 21:{11,11}]
  wire [7:0] _GEN_58 = 8'h3a == io_address ? 8'h3a : _GEN_57; // @[FileReader.scala 21:{11,11}]
  wire [7:0] _GEN_59 = 8'h3b == io_address ? 8'h3b : _GEN_58; // @[FileReader.scala 21:{11,11}]
  wire [7:0] _GEN_60 = 8'h3c == io_address ? 8'h3c : _GEN_59; // @[FileReader.scala 21:{11,11}]
  wire [7:0] _GEN_61 = 8'h3d == io_address ? 8'h3d : _GEN_60; // @[FileReader.scala 21:{11,11}]
  wire [7:0] _GEN_62 = 8'h3e == io_address ? 8'h3e : _GEN_61; // @[FileReader.scala 21:{11,11}]
  wire [7:0] _GEN_63 = 8'h3f == io_address ? 8'h3f : _GEN_62; // @[FileReader.scala 21:{11,11}]
  wire [7:0] _GEN_64 = 8'h40 == io_address ? 8'h40 : _GEN_63; // @[FileReader.scala 21:{11,11}]
  wire [7:0] _GEN_65 = 8'h41 == io_address ? 8'h41 : _GEN_64; // @[FileReader.scala 21:{11,11}]
  wire [7:0] _GEN_66 = 8'h42 == io_address ? 8'h42 : _GEN_65; // @[FileReader.scala 21:{11,11}]
  wire [7:0] _GEN_67 = 8'h43 == io_address ? 8'h43 : _GEN_66; // @[FileReader.scala 21:{11,11}]
  wire [7:0] _GEN_68 = 8'h44 == io_address ? 8'h44 : _GEN_67; // @[FileReader.scala 21:{11,11}]
  wire [7:0] _GEN_69 = 8'h45 == io_address ? 8'h45 : _GEN_68; // @[FileReader.scala 21:{11,11}]
  wire [7:0] _GEN_70 = 8'h46 == io_address ? 8'h46 : _GEN_69; // @[FileReader.scala 21:{11,11}]
  wire [7:0] _GEN_71 = 8'h47 == io_address ? 8'h47 : _GEN_70; // @[FileReader.scala 21:{11,11}]
  wire [7:0] _GEN_72 = 8'h48 == io_address ? 8'h48 : _GEN_71; // @[FileReader.scala 21:{11,11}]
  wire [7:0] _GEN_73 = 8'h49 == io_address ? 8'h49 : _GEN_72; // @[FileReader.scala 21:{11,11}]
  wire [7:0] _GEN_74 = 8'h4a == io_address ? 8'h4a : _GEN_73; // @[FileReader.scala 21:{11,11}]
  wire [7:0] _GEN_75 = 8'h4b == io_address ? 8'h4b : _GEN_74; // @[FileReader.scala 21:{11,11}]
  wire [7:0] _GEN_76 = 8'h4c == io_address ? 8'h4c : _GEN_75; // @[FileReader.scala 21:{11,11}]
  wire [7:0] _GEN_77 = 8'h4d == io_address ? 8'h4d : _GEN_76; // @[FileReader.scala 21:{11,11}]
  wire [7:0] _GEN_78 = 8'h4e == io_address ? 8'h4e : _GEN_77; // @[FileReader.scala 21:{11,11}]
  wire [7:0] _GEN_79 = 8'h4f == io_address ? 8'h4f : _GEN_78; // @[FileReader.scala 21:{11,11}]
  wire [7:0] _GEN_80 = 8'h50 == io_address ? 8'h50 : _GEN_79; // @[FileReader.scala 21:{11,11}]
  wire [7:0] _GEN_81 = 8'h51 == io_address ? 8'h51 : _GEN_80; // @[FileReader.scala 21:{11,11}]
  wire [7:0] _GEN_82 = 8'h52 == io_address ? 8'h52 : _GEN_81; // @[FileReader.scala 21:{11,11}]
  wire [7:0] _GEN_83 = 8'h53 == io_address ? 8'h53 : _GEN_82; // @[FileReader.scala 21:{11,11}]
  wire [7:0] _GEN_84 = 8'h54 == io_address ? 8'h54 : _GEN_83; // @[FileReader.scala 21:{11,11}]
  wire [7:0] _GEN_85 = 8'h55 == io_address ? 8'h55 : _GEN_84; // @[FileReader.scala 21:{11,11}]
  wire [7:0] _GEN_86 = 8'h56 == io_address ? 8'h56 : _GEN_85; // @[FileReader.scala 21:{11,11}]
  wire [7:0] _GEN_87 = 8'h57 == io_address ? 8'h57 : _GEN_86; // @[FileReader.scala 21:{11,11}]
  wire [7:0] _GEN_88 = 8'h58 == io_address ? 8'h58 : _GEN_87; // @[FileReader.scala 21:{11,11}]
  wire [7:0] _GEN_89 = 8'h59 == io_address ? 8'h59 : _GEN_88; // @[FileReader.scala 21:{11,11}]
  wire [7:0] _GEN_90 = 8'h5a == io_address ? 8'h5a : _GEN_89; // @[FileReader.scala 21:{11,11}]
  wire [7:0] _GEN_91 = 8'h5b == io_address ? 8'h5b : _GEN_90; // @[FileReader.scala 21:{11,11}]
  wire [7:0] _GEN_92 = 8'h5c == io_address ? 8'h5c : _GEN_91; // @[FileReader.scala 21:{11,11}]
  wire [7:0] _GEN_93 = 8'h5d == io_address ? 8'h5d : _GEN_92; // @[FileReader.scala 21:{11,11}]
  wire [7:0] _GEN_94 = 8'h5e == io_address ? 8'h5e : _GEN_93; // @[FileReader.scala 21:{11,11}]
  wire [7:0] _GEN_95 = 8'h5f == io_address ? 8'h5f : _GEN_94; // @[FileReader.scala 21:{11,11}]
  wire [7:0] _GEN_96 = 8'h60 == io_address ? 8'h60 : _GEN_95; // @[FileReader.scala 21:{11,11}]
  wire [7:0] _GEN_97 = 8'h61 == io_address ? 8'h61 : _GEN_96; // @[FileReader.scala 21:{11,11}]
  wire [7:0] _GEN_98 = 8'h62 == io_address ? 8'h62 : _GEN_97; // @[FileReader.scala 21:{11,11}]
  wire [7:0] _GEN_99 = 8'h63 == io_address ? 8'h63 : _GEN_98; // @[FileReader.scala 21:{11,11}]
  wire [7:0] _GEN_100 = 8'h64 == io_address ? 8'h64 : _GEN_99; // @[FileReader.scala 21:{11,11}]
  wire [7:0] _GEN_101 = 8'h65 == io_address ? 8'h65 : _GEN_100; // @[FileReader.scala 21:{11,11}]
  wire [7:0] _GEN_102 = 8'h66 == io_address ? 8'h66 : _GEN_101; // @[FileReader.scala 21:{11,11}]
  wire [7:0] _GEN_103 = 8'h67 == io_address ? 8'h67 : _GEN_102; // @[FileReader.scala 21:{11,11}]
  wire [7:0] _GEN_104 = 8'h68 == io_address ? 8'h68 : _GEN_103; // @[FileReader.scala 21:{11,11}]
  wire [7:0] _GEN_105 = 8'h69 == io_address ? 8'h69 : _GEN_104; // @[FileReader.scala 21:{11,11}]
  wire [7:0] _GEN_106 = 8'h6a == io_address ? 8'h6a : _GEN_105; // @[FileReader.scala 21:{11,11}]
  wire [7:0] _GEN_107 = 8'h6b == io_address ? 8'h6b : _GEN_106; // @[FileReader.scala 21:{11,11}]
  wire [7:0] _GEN_108 = 8'h6c == io_address ? 8'h6c : _GEN_107; // @[FileReader.scala 21:{11,11}]
  wire [7:0] _GEN_109 = 8'h6d == io_address ? 8'h6d : _GEN_108; // @[FileReader.scala 21:{11,11}]
  wire [7:0] _GEN_110 = 8'h6e == io_address ? 8'h6e : _GEN_109; // @[FileReader.scala 21:{11,11}]
  wire [7:0] _GEN_111 = 8'h6f == io_address ? 8'h6f : _GEN_110; // @[FileReader.scala 21:{11,11}]
  wire [7:0] _GEN_112 = 8'h70 == io_address ? 8'h70 : _GEN_111; // @[FileReader.scala 21:{11,11}]
  wire [7:0] _GEN_113 = 8'h71 == io_address ? 8'h71 : _GEN_112; // @[FileReader.scala 21:{11,11}]
  wire [7:0] _GEN_114 = 8'h72 == io_address ? 8'h72 : _GEN_113; // @[FileReader.scala 21:{11,11}]
  wire [7:0] _GEN_115 = 8'h73 == io_address ? 8'h73 : _GEN_114; // @[FileReader.scala 21:{11,11}]
  wire [7:0] _GEN_116 = 8'h74 == io_address ? 8'h74 : _GEN_115; // @[FileReader.scala 21:{11,11}]
  wire [7:0] _GEN_117 = 8'h75 == io_address ? 8'h75 : _GEN_116; // @[FileReader.scala 21:{11,11}]
  wire [7:0] _GEN_118 = 8'h76 == io_address ? 8'h76 : _GEN_117; // @[FileReader.scala 21:{11,11}]
  wire [7:0] _GEN_119 = 8'h77 == io_address ? 8'h77 : _GEN_118; // @[FileReader.scala 21:{11,11}]
  wire [7:0] _GEN_120 = 8'h78 == io_address ? 8'h78 : _GEN_119; // @[FileReader.scala 21:{11,11}]
  wire [7:0] _GEN_121 = 8'h79 == io_address ? 8'h79 : _GEN_120; // @[FileReader.scala 21:{11,11}]
  wire [7:0] _GEN_122 = 8'h7a == io_address ? 8'h7a : _GEN_121; // @[FileReader.scala 21:{11,11}]
  wire [7:0] _GEN_123 = 8'h7b == io_address ? 8'h7b : _GEN_122; // @[FileReader.scala 21:{11,11}]
  wire [7:0] _GEN_124 = 8'h7c == io_address ? 8'h7c : _GEN_123; // @[FileReader.scala 21:{11,11}]
  wire [7:0] _GEN_125 = 8'h7d == io_address ? 8'h7d : _GEN_124; // @[FileReader.scala 21:{11,11}]
  wire [7:0] _GEN_126 = 8'h7e == io_address ? 8'h7e : _GEN_125; // @[FileReader.scala 21:{11,11}]
  wire [7:0] _GEN_127 = 8'h7f == io_address ? 8'h7f : _GEN_126; // @[FileReader.scala 21:{11,11}]
  wire [7:0] _GEN_128 = 8'h80 == io_address ? 8'h80 : _GEN_127; // @[FileReader.scala 21:{11,11}]
  wire [7:0] _GEN_129 = 8'h81 == io_address ? 8'h81 : _GEN_128; // @[FileReader.scala 21:{11,11}]
  wire [7:0] _GEN_130 = 8'h82 == io_address ? 8'h82 : _GEN_129; // @[FileReader.scala 21:{11,11}]
  wire [7:0] _GEN_131 = 8'h83 == io_address ? 8'h83 : _GEN_130; // @[FileReader.scala 21:{11,11}]
  wire [7:0] _GEN_132 = 8'h84 == io_address ? 8'h84 : _GEN_131; // @[FileReader.scala 21:{11,11}]
  wire [7:0] _GEN_133 = 8'h85 == io_address ? 8'h85 : _GEN_132; // @[FileReader.scala 21:{11,11}]
  wire [7:0] _GEN_134 = 8'h86 == io_address ? 8'h86 : _GEN_133; // @[FileReader.scala 21:{11,11}]
  wire [7:0] _GEN_135 = 8'h87 == io_address ? 8'h87 : _GEN_134; // @[FileReader.scala 21:{11,11}]
  wire [7:0] _GEN_136 = 8'h88 == io_address ? 8'h88 : _GEN_135; // @[FileReader.scala 21:{11,11}]
  wire [7:0] _GEN_137 = 8'h89 == io_address ? 8'h89 : _GEN_136; // @[FileReader.scala 21:{11,11}]
  wire [7:0] _GEN_138 = 8'h8a == io_address ? 8'h8a : _GEN_137; // @[FileReader.scala 21:{11,11}]
  wire [7:0] _GEN_139 = 8'h8b == io_address ? 8'h8b : _GEN_138; // @[FileReader.scala 21:{11,11}]
  wire [7:0] _GEN_140 = 8'h8c == io_address ? 8'h8c : _GEN_139; // @[FileReader.scala 21:{11,11}]
  wire [7:0] _GEN_141 = 8'h8d == io_address ? 8'h8d : _GEN_140; // @[FileReader.scala 21:{11,11}]
  wire [7:0] _GEN_142 = 8'h8e == io_address ? 8'h8e : _GEN_141; // @[FileReader.scala 21:{11,11}]
  wire [7:0] _GEN_143 = 8'h8f == io_address ? 8'h8f : _GEN_142; // @[FileReader.scala 21:{11,11}]
  wire [7:0] _GEN_144 = 8'h90 == io_address ? 8'h90 : _GEN_143; // @[FileReader.scala 21:{11,11}]
  wire [7:0] _GEN_145 = 8'h91 == io_address ? 8'h91 : _GEN_144; // @[FileReader.scala 21:{11,11}]
  wire [7:0] _GEN_146 = 8'h92 == io_address ? 8'h92 : _GEN_145; // @[FileReader.scala 21:{11,11}]
  wire [7:0] _GEN_147 = 8'h93 == io_address ? 8'h93 : _GEN_146; // @[FileReader.scala 21:{11,11}]
  wire [7:0] _GEN_148 = 8'h94 == io_address ? 8'h94 : _GEN_147; // @[FileReader.scala 21:{11,11}]
  wire [7:0] _GEN_149 = 8'h95 == io_address ? 8'h95 : _GEN_148; // @[FileReader.scala 21:{11,11}]
  wire [7:0] _GEN_150 = 8'h96 == io_address ? 8'h96 : _GEN_149; // @[FileReader.scala 21:{11,11}]
  wire [7:0] _GEN_151 = 8'h97 == io_address ? 8'h97 : _GEN_150; // @[FileReader.scala 21:{11,11}]
  wire [7:0] _GEN_152 = 8'h98 == io_address ? 8'h98 : _GEN_151; // @[FileReader.scala 21:{11,11}]
  wire [7:0] _GEN_153 = 8'h99 == io_address ? 8'h99 : _GEN_152; // @[FileReader.scala 21:{11,11}]
  wire [7:0] _GEN_154 = 8'h9a == io_address ? 8'h9a : _GEN_153; // @[FileReader.scala 21:{11,11}]
  wire [7:0] _GEN_155 = 8'h9b == io_address ? 8'h9b : _GEN_154; // @[FileReader.scala 21:{11,11}]
  wire [7:0] _GEN_156 = 8'h9c == io_address ? 8'h9c : _GEN_155; // @[FileReader.scala 21:{11,11}]
  wire [7:0] _GEN_157 = 8'h9d == io_address ? 8'h9d : _GEN_156; // @[FileReader.scala 21:{11,11}]
  wire [7:0] _GEN_158 = 8'h9e == io_address ? 8'h9e : _GEN_157; // @[FileReader.scala 21:{11,11}]
  wire [7:0] _GEN_159 = 8'h9f == io_address ? 8'h9f : _GEN_158; // @[FileReader.scala 21:{11,11}]
  wire [7:0] _GEN_160 = 8'ha0 == io_address ? 8'ha0 : _GEN_159; // @[FileReader.scala 21:{11,11}]
  wire [7:0] _GEN_161 = 8'ha1 == io_address ? 8'ha1 : _GEN_160; // @[FileReader.scala 21:{11,11}]
  wire [7:0] _GEN_162 = 8'ha2 == io_address ? 8'ha2 : _GEN_161; // @[FileReader.scala 21:{11,11}]
  wire [7:0] _GEN_163 = 8'ha3 == io_address ? 8'ha3 : _GEN_162; // @[FileReader.scala 21:{11,11}]
  wire [7:0] _GEN_164 = 8'ha4 == io_address ? 8'ha4 : _GEN_163; // @[FileReader.scala 21:{11,11}]
  wire [7:0] _GEN_165 = 8'ha5 == io_address ? 8'ha5 : _GEN_164; // @[FileReader.scala 21:{11,11}]
  wire [7:0] _GEN_166 = 8'ha6 == io_address ? 8'ha6 : _GEN_165; // @[FileReader.scala 21:{11,11}]
  wire [7:0] _GEN_167 = 8'ha7 == io_address ? 8'ha7 : _GEN_166; // @[FileReader.scala 21:{11,11}]
  wire [7:0] _GEN_168 = 8'ha8 == io_address ? 8'ha8 : _GEN_167; // @[FileReader.scala 21:{11,11}]
  wire [7:0] _GEN_169 = 8'ha9 == io_address ? 8'ha9 : _GEN_168; // @[FileReader.scala 21:{11,11}]
  wire [7:0] _GEN_170 = 8'haa == io_address ? 8'haa : _GEN_169; // @[FileReader.scala 21:{11,11}]
  wire [7:0] _GEN_171 = 8'hab == io_address ? 8'hab : _GEN_170; // @[FileReader.scala 21:{11,11}]
  wire [7:0] _GEN_172 = 8'hac == io_address ? 8'hac : _GEN_171; // @[FileReader.scala 21:{11,11}]
  wire [7:0] _GEN_173 = 8'had == io_address ? 8'had : _GEN_172; // @[FileReader.scala 21:{11,11}]
  wire [7:0] _GEN_174 = 8'hae == io_address ? 8'hae : _GEN_173; // @[FileReader.scala 21:{11,11}]
  wire [7:0] _GEN_175 = 8'haf == io_address ? 8'haf : _GEN_174; // @[FileReader.scala 21:{11,11}]
  wire [7:0] _GEN_176 = 8'hb0 == io_address ? 8'hb0 : _GEN_175; // @[FileReader.scala 21:{11,11}]
  wire [7:0] _GEN_177 = 8'hb1 == io_address ? 8'hb1 : _GEN_176; // @[FileReader.scala 21:{11,11}]
  wire [7:0] _GEN_178 = 8'hb2 == io_address ? 8'hb2 : _GEN_177; // @[FileReader.scala 21:{11,11}]
  wire [7:0] _GEN_179 = 8'hb3 == io_address ? 8'hb3 : _GEN_178; // @[FileReader.scala 21:{11,11}]
  wire [7:0] _GEN_180 = 8'hb4 == io_address ? 8'hb4 : _GEN_179; // @[FileReader.scala 21:{11,11}]
  wire [7:0] _GEN_181 = 8'hb5 == io_address ? 8'hb5 : _GEN_180; // @[FileReader.scala 21:{11,11}]
  wire [7:0] _GEN_182 = 8'hb6 == io_address ? 8'hb6 : _GEN_181; // @[FileReader.scala 21:{11,11}]
  wire [7:0] _GEN_183 = 8'hb7 == io_address ? 8'hb7 : _GEN_182; // @[FileReader.scala 21:{11,11}]
  wire [7:0] _GEN_184 = 8'hb8 == io_address ? 8'hb8 : _GEN_183; // @[FileReader.scala 21:{11,11}]
  wire [7:0] _GEN_185 = 8'hb9 == io_address ? 8'hb9 : _GEN_184; // @[FileReader.scala 21:{11,11}]
  wire [7:0] _GEN_186 = 8'hba == io_address ? 8'hba : _GEN_185; // @[FileReader.scala 21:{11,11}]
  wire [7:0] _GEN_187 = 8'hbb == io_address ? 8'hbb : _GEN_186; // @[FileReader.scala 21:{11,11}]
  wire [7:0] _GEN_188 = 8'hbc == io_address ? 8'hbc : _GEN_187; // @[FileReader.scala 21:{11,11}]
  wire [7:0] _GEN_189 = 8'hbd == io_address ? 8'hbd : _GEN_188; // @[FileReader.scala 21:{11,11}]
  wire [7:0] _GEN_190 = 8'hbe == io_address ? 8'hbe : _GEN_189; // @[FileReader.scala 21:{11,11}]
  wire [7:0] _GEN_191 = 8'hbf == io_address ? 8'hbf : _GEN_190; // @[FileReader.scala 21:{11,11}]
  wire [7:0] _GEN_192 = 8'hc0 == io_address ? 8'hc0 : _GEN_191; // @[FileReader.scala 21:{11,11}]
  wire [7:0] _GEN_193 = 8'hc1 == io_address ? 8'hc1 : _GEN_192; // @[FileReader.scala 21:{11,11}]
  wire [7:0] _GEN_194 = 8'hc2 == io_address ? 8'hc2 : _GEN_193; // @[FileReader.scala 21:{11,11}]
  wire [7:0] _GEN_195 = 8'hc3 == io_address ? 8'hc3 : _GEN_194; // @[FileReader.scala 21:{11,11}]
  wire [7:0] _GEN_196 = 8'hc4 == io_address ? 8'hc4 : _GEN_195; // @[FileReader.scala 21:{11,11}]
  wire [7:0] _GEN_197 = 8'hc5 == io_address ? 8'hc5 : _GEN_196; // @[FileReader.scala 21:{11,11}]
  wire [7:0] _GEN_198 = 8'hc6 == io_address ? 8'hc6 : _GEN_197; // @[FileReader.scala 21:{11,11}]
  wire [7:0] _GEN_199 = 8'hc7 == io_address ? 8'hc7 : _GEN_198; // @[FileReader.scala 21:{11,11}]
  wire [7:0] _GEN_200 = 8'hc8 == io_address ? 8'hc8 : _GEN_199; // @[FileReader.scala 21:{11,11}]
  wire [7:0] _GEN_201 = 8'hc9 == io_address ? 8'hc9 : _GEN_200; // @[FileReader.scala 21:{11,11}]
  wire [7:0] _GEN_202 = 8'hca == io_address ? 8'hca : _GEN_201; // @[FileReader.scala 21:{11,11}]
  wire [7:0] _GEN_203 = 8'hcb == io_address ? 8'hcb : _GEN_202; // @[FileReader.scala 21:{11,11}]
  wire [7:0] _GEN_204 = 8'hcc == io_address ? 8'hcc : _GEN_203; // @[FileReader.scala 21:{11,11}]
  wire [7:0] _GEN_205 = 8'hcd == io_address ? 8'hcd : _GEN_204; // @[FileReader.scala 21:{11,11}]
  wire [7:0] _GEN_206 = 8'hce == io_address ? 8'hce : _GEN_205; // @[FileReader.scala 21:{11,11}]
  wire [7:0] _GEN_207 = 8'hcf == io_address ? 8'hcf : _GEN_206; // @[FileReader.scala 21:{11,11}]
  wire [7:0] _GEN_208 = 8'hd0 == io_address ? 8'hd0 : _GEN_207; // @[FileReader.scala 21:{11,11}]
  wire [7:0] _GEN_209 = 8'hd1 == io_address ? 8'hd1 : _GEN_208; // @[FileReader.scala 21:{11,11}]
  wire [7:0] _GEN_210 = 8'hd2 == io_address ? 8'hd2 : _GEN_209; // @[FileReader.scala 21:{11,11}]
  wire [7:0] _GEN_211 = 8'hd3 == io_address ? 8'hd3 : _GEN_210; // @[FileReader.scala 21:{11,11}]
  wire [7:0] _GEN_212 = 8'hd4 == io_address ? 8'hd4 : _GEN_211; // @[FileReader.scala 21:{11,11}]
  wire [7:0] _GEN_213 = 8'hd5 == io_address ? 8'hd5 : _GEN_212; // @[FileReader.scala 21:{11,11}]
  wire [7:0] _GEN_214 = 8'hd6 == io_address ? 8'hd6 : _GEN_213; // @[FileReader.scala 21:{11,11}]
  wire [7:0] _GEN_215 = 8'hd7 == io_address ? 8'hd7 : _GEN_214; // @[FileReader.scala 21:{11,11}]
  wire [7:0] _GEN_216 = 8'hd8 == io_address ? 8'hd8 : _GEN_215; // @[FileReader.scala 21:{11,11}]
  wire [7:0] _GEN_217 = 8'hd9 == io_address ? 8'hd9 : _GEN_216; // @[FileReader.scala 21:{11,11}]
  wire [7:0] _GEN_218 = 8'hda == io_address ? 8'hda : _GEN_217; // @[FileReader.scala 21:{11,11}]
  wire [7:0] _GEN_219 = 8'hdb == io_address ? 8'hdb : _GEN_218; // @[FileReader.scala 21:{11,11}]
  wire [7:0] _GEN_220 = 8'hdc == io_address ? 8'hdc : _GEN_219; // @[FileReader.scala 21:{11,11}]
  wire [7:0] _GEN_221 = 8'hdd == io_address ? 8'hdd : _GEN_220; // @[FileReader.scala 21:{11,11}]
  wire [7:0] _GEN_222 = 8'hde == io_address ? 8'hde : _GEN_221; // @[FileReader.scala 21:{11,11}]
  wire [7:0] _GEN_223 = 8'hdf == io_address ? 8'hdf : _GEN_222; // @[FileReader.scala 21:{11,11}]
  wire [7:0] _GEN_224 = 8'he0 == io_address ? 8'he0 : _GEN_223; // @[FileReader.scala 21:{11,11}]
  wire [7:0] _GEN_225 = 8'he1 == io_address ? 8'he1 : _GEN_224; // @[FileReader.scala 21:{11,11}]
  wire [7:0] _GEN_226 = 8'he2 == io_address ? 8'he2 : _GEN_225; // @[FileReader.scala 21:{11,11}]
  wire [7:0] _GEN_227 = 8'he3 == io_address ? 8'he3 : _GEN_226; // @[FileReader.scala 21:{11,11}]
  wire [7:0] _GEN_228 = 8'he4 == io_address ? 8'he4 : _GEN_227; // @[FileReader.scala 21:{11,11}]
  wire [7:0] _GEN_229 = 8'he5 == io_address ? 8'he5 : _GEN_228; // @[FileReader.scala 21:{11,11}]
  wire [7:0] _GEN_230 = 8'he6 == io_address ? 8'he6 : _GEN_229; // @[FileReader.scala 21:{11,11}]
  wire [7:0] _GEN_231 = 8'he7 == io_address ? 8'he7 : _GEN_230; // @[FileReader.scala 21:{11,11}]
  wire [7:0] _GEN_232 = 8'he8 == io_address ? 8'he8 : _GEN_231; // @[FileReader.scala 21:{11,11}]
  wire [7:0] _GEN_233 = 8'he9 == io_address ? 8'he9 : _GEN_232; // @[FileReader.scala 21:{11,11}]
  wire [7:0] _GEN_234 = 8'hea == io_address ? 8'hea : _GEN_233; // @[FileReader.scala 21:{11,11}]
  wire [7:0] _GEN_235 = 8'heb == io_address ? 8'heb : _GEN_234; // @[FileReader.scala 21:{11,11}]
  wire [7:0] _GEN_236 = 8'hec == io_address ? 8'hec : _GEN_235; // @[FileReader.scala 21:{11,11}]
  wire [7:0] _GEN_237 = 8'hed == io_address ? 8'hed : _GEN_236; // @[FileReader.scala 21:{11,11}]
  wire [7:0] _GEN_238 = 8'hee == io_address ? 8'hee : _GEN_237; // @[FileReader.scala 21:{11,11}]
  wire [7:0] _GEN_239 = 8'hef == io_address ? 8'hef : _GEN_238; // @[FileReader.scala 21:{11,11}]
  wire [7:0] _GEN_240 = 8'hf0 == io_address ? 8'hf0 : _GEN_239; // @[FileReader.scala 21:{11,11}]
  wire [7:0] _GEN_241 = 8'hf1 == io_address ? 8'hf1 : _GEN_240; // @[FileReader.scala 21:{11,11}]
  wire [7:0] _GEN_242 = 8'hf2 == io_address ? 8'hf2 : _GEN_241; // @[FileReader.scala 21:{11,11}]
  wire [7:0] _GEN_243 = 8'hf3 == io_address ? 8'hf3 : _GEN_242; // @[FileReader.scala 21:{11,11}]
  wire [7:0] _GEN_244 = 8'hf4 == io_address ? 8'hf4 : _GEN_243; // @[FileReader.scala 21:{11,11}]
  wire [7:0] _GEN_245 = 8'hf5 == io_address ? 8'hf5 : _GEN_244; // @[FileReader.scala 21:{11,11}]
  wire [7:0] _GEN_246 = 8'hf6 == io_address ? 8'hf6 : _GEN_245; // @[FileReader.scala 21:{11,11}]
  wire [7:0] _GEN_247 = 8'hf7 == io_address ? 8'hf7 : _GEN_246; // @[FileReader.scala 21:{11,11}]
  wire [7:0] _GEN_248 = 8'hf8 == io_address ? 8'hf8 : _GEN_247; // @[FileReader.scala 21:{11,11}]
  wire [7:0] _GEN_249 = 8'hf9 == io_address ? 8'hf9 : _GEN_248; // @[FileReader.scala 21:{11,11}]
  wire [7:0] _GEN_250 = 8'hfa == io_address ? 8'hfa : _GEN_249; // @[FileReader.scala 21:{11,11}]
  wire [7:0] _GEN_251 = 8'hfb == io_address ? 8'hfb : _GEN_250; // @[FileReader.scala 21:{11,11}]
  wire [7:0] _GEN_252 = 8'hfc == io_address ? 8'hfc : _GEN_251; // @[FileReader.scala 21:{11,11}]
  wire [7:0] _GEN_253 = 8'hfd == io_address ? 8'hfd : _GEN_252; // @[FileReader.scala 21:{11,11}]
  wire [7:0] _GEN_254 = 8'hfe == io_address ? 8'hfe : _GEN_253; // @[FileReader.scala 21:{11,11}]
  assign io_data = 8'hff == io_address ? 8'hff : _GEN_254; // @[FileReader.scala 21:{11,11}]
endmodule
